//  ************    CFLib   *******************************************
//
//  Organisation:   Chipforge
//                  Germany / European Union
//
//  Profile:        Chipforge focus on fine System-on-Chip Cores in
//                  Verilog HDL Code which are easy understandable and
//                  adjustable. For further information see
//                          www.chipforge.org
//                  there are projects from small cores up to PCBs, too.
//
//  File:           CFLib/asyncrst/TBench/tb_asyncrst.sv
//
//  Purpose:        Test Bench for asyncrst
//
//  ************    IEEE 1800-2012 (SystemVerilog 2012) ***************
//
//  ///////////////////////////////////////////////////////////////////
//
//  Copyright (c)   2019, 2020 by
//                  chipforge <cflib@nospam.chipforge.org>
//
//      This Source Code Library is licensed under the Libre Silicon
//      public license; you can redistribute it and/or modify it under
//      the terms of the Libre Silicon public license as published by
//      the Libre Silicon alliance, either version 1 of the License, or
//      (at your option) any later version.
//
//      This design is distributed in the hope that it will be useful,
//      but WITHOUT ANY WARRANTY; without even the implied warranty of
//      MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.
//      See the Libre Silicon Public License for more details.
//
//  ///////////////////////////////////////////////////////////////////

